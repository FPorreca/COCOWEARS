constant A_MATRIX : COEFF_MATRIX := (
    0 => (
        "000000000000100000000000000000"  --(1.000000000000),
        "111111111111011000110101111000"  --(-1.223693847656),
        "000000000000001101111011101010"  --(0.435379028320)
    ),
    1 => (
        "000000000000100000000000000000"  --(1.000000000000),
        "111111111111010110111010111000"  --(-1.283752441406),
        "000000000000010110100000100111"  --(0.703422546387)
    ),
    2 => (
        "000000000000100000000000000000"  --(1.000000000000),
        "111111111111001001011110110010"  --(-1.703720092773),
        "000000000000010111101000111011"  --(0.738731384277)
    ),
    3 => (
        "000000000000100000000000000000"  --(1.000000000000),
        "111111111111000011001010101000"  --(-1.901062011719),
        "000000000000011101100010100001"  --(0.923103332520)
    )
);

constant B_MATRIX : COEFF_MATRIX := (
    0 => (
        "000000000000000000000111111011"  --(0.003868103027),
        "000000000000000000001111110110"  --(0.007736206055),
        "000000000000000000000111111011"  --(0.003868103027)
    ),
    1 => (
        "000000000000100000000000000000"  --(1.000000000000),
        "000000000001000000000000000000"  --(2.000000000000),
        "000000000000100000000000000000"  --(1.000000000000)
    ),
    2 => (
        "000000000000100000000000000000"  --(1.000000000000),
        "111111111111000000000000000000"  --(-2.000000000000),
        "000000000000100000000000000000"  --(1.000000000000)
    ),
    3 => (
        "000000000000100000000000000000"  --(1.000000000000),
        "111111111111000000000000000000"  --(-2.000000000000),
        "000000000000100000000000000000"  --(1.000000000000)
    )
);
