library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity testbench is
end entity testbench;

architecture sim of testbench is
    component iir_filter
        port (
            clk : in  std_logic;
            rst : in  std_logic;
            x   : in  std_logic_vector(17 downto 0);
            y   : out std_logic_vector(17 downto 0)
        );
    end component;

    signal clk : std_logic := '0';
    signal rst : std_logic := '1';
    signal x   : std_logic_vector(17 downto 0) := (others => '0');
    signal y   : std_logic_vector(17 downto 0);

    constant clk_period : time := 11.6 ns;
    constant start_time : time := 360 ns;
    constant stop_time : time := 11960 ns;
begin

    
    clk_process : process
    begin
        while true loop
            clk <= '0';
            wait for clk_period / 2;
            clk <= '1';
            wait for clk_period / 2;
        end loop;
    end process;

    
    uut: iir_filter
        port map (
            clk => clk,
            rst => rst,
            x   => x,
            y   => y
        );

    
    stim_proc : process
        begin
            wait for 102ns;
            rst <= '0';
x <= "111111110111111010";  
wait for clk_period;
x <= "000001101011101111";  
wait for clk_period;
x <= "000010000011001111";  
wait for clk_period;
x <= "000000111111110110";  
wait for clk_period;
x <= "000000000100110100";  
wait for clk_period;
x <= "111111110010101000";  
wait for clk_period;
x <= "111111110101110011";  
wait for clk_period;
x <= "000000100001001010";  
wait for clk_period;
x <= "000000101001001000";  
wait for clk_period;
x <= "000001001101001101";  
wait for clk_period;
x <= "000000100001110001";  
wait for clk_period;
x <= "000010000101010001";  
wait for clk_period;
x <= "111110110000101111";  
wait for clk_period;
x <= "111111110000111101";  
wait for clk_period;
x <= "111111001000000110";  
wait for clk_period;
x <= "000000111011000100";  
wait for clk_period;
x <= "111111100010110000";  
wait for clk_period;
x <= "111111100000100111";  
wait for clk_period;
x <= "000001111101011010";  
wait for clk_period;
x <= "000000001001100010";  
wait for clk_period;
x <= "000000011100101011";  
wait for clk_period;
x <= "111111010010111010";  
wait for clk_period;
x <= "000001001101100011";  
wait for clk_period;
x <= "111111011011110110";  
wait for clk_period;
x <= "000000010101000010";  
wait for clk_period;
x <= "111111110111111101";  
wait for clk_period;
x <= "000000001010000011";  
wait for clk_period;
x <= "000000111010010100";  
wait for clk_period;
x <= "000000111100100100";  
wait for clk_period;
x <= "111110001110001001";  
wait for clk_period;
x <= "000000000101010010";  
wait for clk_period;
x <= "111111111010111100";  
wait for clk_period;
x <= "111111001011001011";  
wait for clk_period;
x <= "111111000100110110";  
wait for clk_period;
x <= "111110110011101000";  
wait for clk_period;
x <= "000000000111110010";  
wait for clk_period;
x <= "000000010000101110";  
wait for clk_period;
x <= "000001101010100100";  
wait for clk_period;
x <= "111110101000100000";  
wait for clk_period;
x <= "000000000110001101";  
wait for clk_period;
x <= "111101110010001010";  
wait for clk_period;
x <= "111110010101001010";  
wait for clk_period;
x <= "000000111001001001";  
wait for clk_period;
x <= "000000101000001000";  
wait for clk_period;
x <= "000000001110000110";  
wait for clk_period;
x <= "000001000000110011";  
wait for clk_period;
x <= "111111000101000110";  
wait for clk_period;
x <= "111101110000010100";  
wait for clk_period;
x <= "111111100001001101";  
wait for clk_period;
x <= "000000101000100101";  
wait for clk_period;
x <= "111111110101110000";  
wait for clk_period;
x <= "000001010011101011";  
wait for clk_period;
x <= "000001010111101000";  
wait for clk_period;
x <= "000000001111101100";  
wait for clk_period;
x <= "000000001110101101";  
wait for clk_period;
x <= "111111000000010110";  
wait for clk_period;
x <= "000000001011000100";  
wait for clk_period;
x <= "000000011110000101";  
wait for clk_period;
x <= "000000101000110000";  
wait for clk_period;
x <= "111111100111010011";  
wait for clk_period;
x <= "000000100001100111";  
wait for clk_period;
x <= "111111000000110000";  
wait for clk_period;
x <= "000000100001001111";  
wait for clk_period;
x <= "111110101110100100";  
wait for clk_period;
x <= "111111010101100001";  
wait for clk_period;
x <= "111111111010001110";  
wait for clk_period;
x <= "111111100010000110";  
wait for clk_period;
x <= "000000010100011110";  
wait for clk_period;
x <= "111111111000000010";  
wait for clk_period;
x <= "000001101011010111";  
wait for clk_period;
x <= "111111000100111011";  
wait for clk_period;
x <= "000000011100001100";  
wait for clk_period;
x <= "000000001010110010";  
wait for clk_period;
x <= "000001101111110111";  
wait for clk_period;
x <= "000000000100111001";  
wait for clk_period;
x <= "111111000001110101";  
wait for clk_period;
x <= "000000001111110010";  
wait for clk_period;
x <= "000000111111000111";  
wait for clk_period;
x <= "111111100101110111";  
wait for clk_period;
x <= "111111111000101110";  
wait for clk_period;
x <= "000000000010100011";  
wait for clk_period;
x <= "111111011001100101";  
wait for clk_period;
x <= "111110110010101001";  
wait for clk_period;
x <= "111110101110010100";  
wait for clk_period;
x <= "000000001100101100";  
wait for clk_period;
x <= "000000011011101000";  
wait for clk_period;
x <= "000001111001100010";  
wait for clk_period;
x <= "111110111011111101";  
wait for clk_period;
x <= "000000001010101011";  
wait for clk_period;
x <= "000000010110110101";  
wait for clk_period;
x <= "000000100001111011";  
wait for clk_period;
x <= "111111110010100001";  
wait for clk_period;
x <= "000000110100011000";  
wait for clk_period;
x <= "000010110000001110";  
wait for clk_period;
x <= "000000101011001011";  
wait for clk_period;
x <= "111111001111001110";  
wait for clk_period;
x <= "111111001111011110";  
wait for clk_period;
x <= "111111100100110111";  
wait for clk_period;
x <= "000000111000010010";  
wait for clk_period;
x <= "000000011100100101";  
wait for clk_period;
x <= "111111110001011101";  
wait for clk_period;
x <= "111111101001110011";  
wait for clk_period;
x <= "000000000000100010";  
wait for clk_period;
x <= "000000000000001010";  
wait for clk_period;
x <= "111110111011010110";  
wait for clk_period;
x <= "111111111110111001";  
wait for clk_period;
x <= "111110111101100000";  
wait for clk_period;
x <= "000001001101001000";  
wait for clk_period;
x <= "111111110100110111";  
wait for clk_period;
x <= "111111100001010111";  
wait for clk_period;
x <= "111111110111001000";  
wait for clk_period;
x <= "000000011001011101";  
wait for clk_period;
x <= "111101111010000011";  
wait for clk_period;
x <= "111111000000100101";  
wait for clk_period;
x <= "000000101100010011";  
wait for clk_period;
x <= "111111011110011111";  
wait for clk_period;
x <= "000000100010011010";  
wait for clk_period;
x <= "111110100011110000";  
wait for clk_period;
x <= "111111001000110100";  
wait for clk_period;
x <= "111111110110011101";  
wait for clk_period;
x <= "000001000011011110";  
wait for clk_period;
x <= "111110010101110000";  
wait for clk_period;
x <= "000000000010101110";  
wait for clk_period;
x <= "000000111000000100";  
wait for clk_period;
x <= "111111110010011000";  
wait for clk_period;
x <= "111111110010000001";  
wait for clk_period;
x <= "111110110001111111";  
wait for clk_period;
x <= "000000011010101110";  
wait for clk_period;
x <= "000001000100010101";  
wait for clk_period;
x <= "111111011011110111";  
wait for clk_period;
x <= "111111000100000011";  
wait for clk_period;
x <= "111111111100000010";  
wait for clk_period;
x <= "111111101101000111";  
wait for clk_period;
x <= "000000000111001001";  
wait for clk_period;
x <= "000001000011011001";  
wait for clk_period;
x <= "000010000000110011";  
wait for clk_period;
x <= "111111101010101100";  
wait for clk_period;
x <= "000000001101110110";  
wait for clk_period;
x <= "111111100000111111";  
wait for clk_period;
x <= "000001001001111101";  
wait for clk_period;
x <= "000010001010110011";  
wait for clk_period;
x <= "000001001001001111";  
wait for clk_period;
x <= "000001010100011111";  
wait for clk_period;
x <= "000000011111110011";  
wait for clk_period;
x <= "111111111111011111";  
wait for clk_period;
x <= "111111111110011011";  
wait for clk_period;
x <= "111111000010111011";  
wait for clk_period;
x <= "000000001001101101";  
wait for clk_period;
x <= "000000100110010100";  
wait for clk_period;
x <= "000000000101101101";  
wait for clk_period;
x <= "111111111011000100";  
wait for clk_period;
x <= "000000100110110111";  
wait for clk_period;
x <= "111111100010111101";  
wait for clk_period;
x <= "111101010001101010";  
wait for clk_period;
x <= "000000011101001010";  
wait for clk_period;
x <= "111111101010001100";  
wait for clk_period;
x <= "000001000001010011";  
wait for clk_period;
x <= "000000011101100001";  
wait for clk_period;
x <= "000000101100010000";  
wait for clk_period;
x <= "000000001101101100";  
wait for clk_period;
x <= "111111110010000001";  
wait for clk_period;
x <= "111111101001111001";  
wait for clk_period;
x <= "111110100000011011";  
wait for clk_period;
x <= "000000011100000100";  
wait for clk_period;
x <= "000000000100000001";  
wait for clk_period;
x <= "000000110101100100";  
wait for clk_period;
x <= "111110110101100110";  
wait for clk_period;
x <= "111110111110011111";  
wait for clk_period;
x <= "111110010011110000";  
wait for clk_period;
x <= "000000000011110010";  
wait for clk_period;
x <= "111111011011010111";  
wait for clk_period;
x <= "111111000110010111";  
wait for clk_period;
x <= "111111110100111101";  
wait for clk_period;
x <= "111111100011111010";  
wait for clk_period;
x <= "000000000100001010";  
wait for clk_period;
x <= "000000000111101100";  
wait for clk_period;
x <= "000001001101011001";  
wait for clk_period;
x <= "000000000001011110";  
wait for clk_period;
x <= "111111110010111010";  
wait for clk_period;
x <= "111111101101001000";  
wait for clk_period;
x <= "111110011110011001";  
wait for clk_period;
x <= "000001001010001011";  
wait for clk_period;
x <= "000010001000101001";  
wait for clk_period;
x <= "111111100011111111";  
wait for clk_period;
x <= "000000000001011010";  
wait for clk_period;
x <= "000000110001000110";  
wait for clk_period;
x <= "000000001100001010";  
wait for clk_period;
x <= "111110001110000110";  
wait for clk_period;
x <= "111111101001011000";  
wait for clk_period;
x <= "000000010101011111";  
wait for clk_period;
x <= "000001100000101101";  
wait for clk_period;
x <= "000001101100110011";  
wait for clk_period;
x <= "111111011001011011";  
wait for clk_period;
x <= "000000011010000001";  
wait for clk_period;
x <= "111111111110001010";  
wait for clk_period;
x <= "111110110000001011";  
wait for clk_period;
x <= "111111111101101001";  
wait for clk_period;
x <= "000000000110010010";  
wait for clk_period;
x <= "000000010101100111";  
wait for clk_period;
x <= "000001000011011110";  
wait for clk_period;
x <= "000000010110111011";  
wait for clk_period;
x <= "111111101111000011";  
wait for clk_period;
x <= "111110111000101101";  
wait for clk_period;
x <= "111111111101100101";  
wait for clk_period;
x <= "111110011100011111";  
wait for clk_period;
x <= "000001001011001100";  
wait for clk_period;
x <= "000001100100000011";  
wait for clk_period;
x <= "000000101100111011";  
wait for clk_period;
x <= "000000110111111110";  
wait for clk_period;
x <= "111111100110001110";  
wait for clk_period;
x <= "111111110100000111";  
wait for clk_period;
x <= "111110111101101100";  
wait for clk_period;
x <= "000000101000011011";  
wait for clk_period;
x <= "000000001101110010";  
wait for clk_period;
x <= "111111110001111110";  
wait for clk_period;
x <= "111111000100111100";  
wait for clk_period;
x <= "000000101111010101";  
wait for clk_period;
x <= "000000100110010001";  
wait for clk_period;
x <= "111111000100010111";  
wait for clk_period;
x <= "111111100010101111";  
wait for clk_period;
x <= "111111100111000001";  
wait for clk_period;
x <= "111111101111011011";  
wait for clk_period;
x <= "111111110110111111";  
wait for clk_period;
x <= "000000111100000001";  
wait for clk_period;
x <= "000000010110011100";  
wait for clk_period;
x <= "000001111111011000";  
wait for clk_period;
x <= "000001010001111101";  
wait for clk_period;
x <= "111111010001110111";  
wait for clk_period;
x <= "111111101010000000";  
wait for clk_period;
x <= "111111001111110000";  
wait for clk_period;
x <= "111111111101101111";  
wait for clk_period;
x <= "000000010101111110";  
wait for clk_period;
x <= "000000111100110011";  
wait for clk_period;
x <= "000000010010001100";  
wait for clk_period;
x <= "111111001011100110";  
wait for clk_period;
x <= "111110110101110011";  
wait for clk_period;
x <= "111110000011110100";  
wait for clk_period;
x <= "111111111010000000";  
wait for clk_period;
x <= "111110101110111110";  
wait for clk_period;
x <= "111111000110111101";  
wait for clk_period;
x <= "000000111011000110";  
wait for clk_period;
x <= "000000001010111110";  
wait for clk_period;
x <= "000000001100000000";  
wait for clk_period;
x <= "000000000110110101";  
wait for clk_period;
x <= "111111001001001010";  
wait for clk_period;
x <= "111110010101111110";  
wait for clk_period;
x <= "111111000000010010";  
wait for clk_period;
x <= "000001100101101010";  
wait for clk_period;
x <= "000000101001101011";  
wait for clk_period;
x <= "111111110101110000";  
wait for clk_period;
x <= "000000011111011001";  
wait for clk_period;
x <= "111110110100011101";  
wait for clk_period;
x <= "111111011111101100";  
wait for clk_period;
x <= "111111000000000100";  
wait for clk_period;
x <= "000000001100110011";  
wait for clk_period;
x <= "111111101011001101";  
wait for clk_period;
x <= "000001000010110100";  
wait for clk_period;
x <= "000000101101000111";  
wait for clk_period;
x <= "111111001001001101";  
wait for clk_period;
x <= "000001001100101111";  
wait for clk_period;
x <= "111111100011010110";  
wait for clk_period;
x <= "000000010100001001";  
wait for clk_period;
x <= "000000100001101011";  
wait for clk_period;
x <= "000000001101101100";  
wait for clk_period;
x <= "000000100100111111";  
wait for clk_period;
x <= "000000011010000101";  
wait for clk_period;
x <= "000001001010010010";  
wait for clk_period;
x <= "000000101111111000";  
wait for clk_period;
x <= "000001110111000110";  
wait for clk_period;
x <= "111110100100001011";  
wait for clk_period;
x <= "111111011110010010";  
wait for clk_period;
x <= "000001000100010000";  
wait for clk_period;
x <= "000000001100110111";  
wait for clk_period;
x <= "000000100111000011";  
wait for clk_period;
x <= "000001110000001001";  
wait for clk_period;
x <= "000000110011111100";  
wait for clk_period;
x <= "111111000101011110";  
wait for clk_period;
x <= "000000000110010111";  
wait for clk_period;
x <= "111111100111110100";  
wait for clk_period;
x <= "000000100010100010";  
wait for clk_period;
x <= "111111011101110001";  
wait for clk_period;
x <= "111111010010111010";  
wait for clk_period;
x <= "000000011001011100";  
wait for clk_period;
x <= "000000011010000001";  
wait for clk_period;
x <= "111111100101001010";  
wait for clk_period;
x <= "111101111100111101";  
wait for clk_period;
x <= "111110101101111110";  
wait for clk_period;
x <= "111111010110000011";  
wait for clk_period;
x <= "000000011110000110";  
wait for clk_period;
x <= "111111001100010001";  
wait for clk_period;
x <= "111111101100000111";  
wait for clk_period;
x <= "000001100010010000";  
wait for clk_period;
x <= "111111110011011010";  
wait for clk_period;
x <= "111110111011011110";  
wait for clk_period;
x <= "111111100100000101";  
wait for clk_period;
x <= "111111110001110001";  
wait for clk_period;
x <= "000000110110011000";  
wait for clk_period;
x <= "000000010000111101";  
wait for clk_period;
x <= "000000000001111110";  
wait for clk_period;
x <= "111111111110010101";  
wait for clk_period;
x <= "111111100111000110";  
wait for clk_period;
x <= "111110100100111001";  
wait for clk_period;
x <= "111110111101101011";  
wait for clk_period;
x <= "000000010001111000";  
wait for clk_period;
x <= "111111100000100010";  
wait for clk_period;
x <= "000000011001111101";  
wait for clk_period;
x <= "111111100010111111";  
wait for clk_period;
x <= "111110100000101110";  
wait for clk_period;
x <= "000001100100111011";  
wait for clk_period;
x <= "000001000111010110";  
wait for clk_period;
x <= "111111111010011010";  
wait for clk_period;
x <= "111111111110000001";  
wait for clk_period;
x <= "000000101101011001";  
wait for clk_period;
x <= "000001011110101010";  
wait for clk_period;
x <= "000000011110000010";  
wait for clk_period;
x <= "000001010101101111";  
wait for clk_period;
x <= "111111010000101111";  
wait for clk_period;
x <= "000000111111010001";  
wait for clk_period;
x <= "000000011011110000";  
wait for clk_period;
x <= "111111000011011000";  
wait for clk_period;
x <= "111111101001110000";  
wait for clk_period;
x <= "000000001100000111";  
wait for clk_period;
x <= "000000111010010100";  
wait for clk_period;
x <= "111110110110101001";  
wait for clk_period;
x <= "111111110101110010";  
wait for clk_period;
x <= "111111111101110100";  
wait for clk_period;
x <= "000000011100100000";  
wait for clk_period;
x <= "111110111110001100";  
wait for clk_period;
x <= "111111110010011100";  
wait for clk_period;
x <= "000000110010110100";  
wait for clk_period;
x <= "000000110110111001";  
wait for clk_period;
x <= "111111010101111001";  
wait for clk_period;
x <= "111111011000111100";  
wait for clk_period;
x <= "000001001010100010";  
wait for clk_period;
x <= "111111111101001110";  
wait for clk_period;
x <= "111111100001111000";  
wait for clk_period;
x <= "111111100100001000";  
wait for clk_period;
x <= "000000010001110111";  
wait for clk_period;
x <= "000000010010010000";  
wait for clk_period;
x <= "000000110000101010";  
wait for clk_period;
x <= "000000001110001101";  
wait for clk_period;
x <= "111110111010011011";  
wait for clk_period;
x <= "111111111111001000";  
wait for clk_period;
x <= "111111011000111010";  
wait for clk_period;
x <= "111111100100001000";  
wait for clk_period;
x <= "000010000101101011";  
wait for clk_period;
x <= "000000100001101010";  
wait for clk_period;
x <= "111111101100111011";  
wait for clk_period;
x <= "111111001111101010";  
wait for clk_period;
x <= "000000001111011111";  
wait for clk_period;
x <= "111111111001111110";  
wait for clk_period;
x <= "111111001111110001";  
wait for clk_period;
x <= "111111101100101110";  
wait for clk_period;
x <= "000000000101010011";  
wait for clk_period;
x <= "000000110010101111";  
wait for clk_period;
x <= "111111100101110101";  
wait for clk_period;
x <= "000000000001100100";  
wait for clk_period;
x <= "000000011111100111";  
wait for clk_period;
x <= "111111101110100001";  
wait for clk_period;
x <= "111111111101011001";  
wait for clk_period;
x <= "000000010101111011";  
wait for clk_period;
x <= "111111100000101111";  
wait for clk_period;
x <= "000001110010010100";  
wait for clk_period;
x <= "111111110100111001";  
wait for clk_period;
x <= "000000100011011001";  
wait for clk_period;
x <= "111111000011000101";  
wait for clk_period;
x <= "111111011000000011";  
wait for clk_period;
x <= "111110101101110110";  
wait for clk_period;
x <= "111110101111111101";  
wait for clk_period;
x <= "111111101000000110";  
wait for clk_period;
x <= "111111011111100110";  
wait for clk_period;
x <= "000001101110000111";  
wait for clk_period;
x <= "111101111010101000";  
wait for clk_period;
x <= "111111000011101100";  
wait for clk_period;
x <= "111111011001010011";  
wait for clk_period;
x <= "111111110101101101";  
wait for clk_period;
x <= "111111110000001000";  
wait for clk_period;
x <= "000000011011011100";  
wait for clk_period;
x <= "111111011101000011";  
wait for clk_period;
x <= "000001001100010101";  
wait for clk_period;
x <= "000010011011110011";  
wait for clk_period;
x <= "111111111010011110";  
wait for clk_period;
x <= "111111010110000110";  
wait for clk_period;
x <= "000000110000110110";  
wait for clk_period;
x <= "111111110010100111";  
wait for clk_period;
x <= "111111010001100111";  
wait for clk_period;
x <= "000000101010001010";  
wait for clk_period;
x <= "000000110100101000";  
wait for clk_period;
x <= "000001001011000100";  
wait for clk_period;
x <= "000000000011010000";  
wait for clk_period;
x <= "111110011011010010";  
wait for clk_period;
x <= "111111101111011100";  
wait for clk_period;
x <= "000000100010001111";  
wait for clk_period;
x <= "111111010110011101";  
wait for clk_period;
x <= "000000111011011101";  
wait for clk_period;
x <= "000000111011100111";  
wait for clk_period;
x <= "000001101110111010";  
wait for clk_period;
x <= "000000100100010010";  
wait for clk_period;
x <= "000000011010101011";  
wait for clk_period;
x <= "111111011101101101";  
wait for clk_period;
x <= "000000110010100000";  
wait for clk_period;
x <= "000001000101101100";  
wait for clk_period;
x <= "111111011000110101";  
wait for clk_period;
x <= "000000100000101101";  
wait for clk_period;
x <= "000001000011111100";  
wait for clk_period;
x <= "000001010110101010";  
wait for clk_period;
x <= "111111011011000011";  
wait for clk_period;
x <= "111111101000101001";  
wait for clk_period;
x <= "111110101100111010";  
wait for clk_period;
x <= "111110101000000001";  
wait for clk_period;
x <= "111111010011100001";  
wait for clk_period;
x <= "000001101100100101";  
wait for clk_period;
x <= "111111100110000010";  
wait for clk_period;
x <= "000000000011110010";  
wait for clk_period;
x <= "111111000110101110";  
wait for clk_period;
x <= "111111000010011000";  
wait for clk_period;
x <= "111110101111011011";  
wait for clk_period;
x <= "111110110011100101";  
wait for clk_period;
x <= "000000010100011001";  
wait for clk_period;
x <= "111110111101101000";  
wait for clk_period;
x <= "000001001010000111";  
wait for clk_period;
x <= "111110101010111010";  
wait for clk_period;
x <= "000000101011111101";  
wait for clk_period;
x <= "111111001100010110";  
wait for clk_period;
x <= "111111000000010001";  
wait for clk_period;
x <= "111111001100010011";  
wait for clk_period;
x <= "111111000010110010";  
wait for clk_period;
x <= "000000100001000100";  
wait for clk_period;
x <= "000000100101110100";  
wait for clk_period;
x <= "000000101100110101";  
wait for clk_period;
x <= "000000011111101011";  
wait for clk_period;
x <= "000000101001101101";  
wait for clk_period;
x <= "111111101011011000";  
wait for clk_period;
x <= "111110100100001111";  
wait for clk_period;
x <= "111111010110110001";  
wait for clk_period;
x <= "000000011111100011";  
wait for clk_period;
x <= "000000100110111100";  
wait for clk_period;
x <= "000000111110000000";  
wait for clk_period;
x <= "111111110100001001";  
wait for clk_period;
x <= "000000000110000010";  
wait for clk_period;
x <= "111110111010111101";  
wait for clk_period;
x <= "111111111001000101";  
wait for clk_period;
x <= "000000011010111101";  
wait for clk_period;
x <= "000000000010100101";  
wait for clk_period;
x <= "111111011111001111";  
wait for clk_period;
x <= "000010011111001101";  
wait for clk_period;
x <= "000001000110101001";  
wait for clk_period;
x <= "000000111011110001";  
wait for clk_period;
x <= "000001000011111110";  
wait for clk_period;
x <= "111111101100001001";  
wait for clk_period;
x <= "111111100010001101";  
wait for clk_period;
x <= "111111110001011001";  
wait for clk_period;
x <= "000000110010000101";  
wait for clk_period;
x <= "111111101111100011";  
wait for clk_period;
x <= "000010000010001010";  
wait for clk_period;
x <= "111110101111010100";  
wait for clk_period;
x <= "111110110001100000";  
wait for clk_period;
x <= "111111011000000001";  
wait for clk_period;
x <= "111111001000110111";  
wait for clk_period;
x <= "111110101011101100";  
wait for clk_period;
x <= "000000011001010001";  
wait for clk_period;
x <= "111111101111111011";  
wait for clk_period;
x <= "000001101001100000";  
wait for clk_period;
x <= "000000110101000100";  
wait for clk_period;
x <= "111111001001111111";  
wait for clk_period;
x <= "111111101111001011";  
wait for clk_period;
x <= "000000001001101111";  
wait for clk_period;
x <= "000000010010011011";  
wait for clk_period;
x <= "111110111011100110";  
wait for clk_period;
x <= "000001111101001110";  
wait for clk_period;
x <= "111110111111010010";  
wait for clk_period;
x <= "000000100110010101";  
wait for clk_period;
x <= "000000101110000100";  
wait for clk_period;
x <= "000000001000110100";  
wait for clk_period;
x <= "111110101101110011";  
wait for clk_period;
x <= "111110011100100110";  
wait for clk_period;
x <= "000000001001110110";  
wait for clk_period;
x <= "000000001000111100";  
wait for clk_period;
x <= "000000110011000110";  
wait for clk_period;
x <= "111111111100101101";  
wait for clk_period;
x <= "111111100101001001";  
wait for clk_period;
x <= "000000001100110111";  
wait for clk_period;
x <= "111111100100111010";  
wait for clk_period;
x <= "111111100000101001";  
wait for clk_period;
x <= "111111111001010010";  
wait for clk_period;
x <= "000000100100101001";  
wait for clk_period;
x <= "000000100010100100";  
wait for clk_period;
x <= "111111000111010001";  
wait for clk_period;
x <= "000000110111001111";  
wait for clk_period;
x <= "000000001110010110";  
wait for clk_period;
x <= "000000010100001110";  
wait for clk_period;
x <= "111110000001101001";  
wait for clk_period;
x <= "111111010001101100";  
wait for clk_period;
x <= "111111111010100100";  
wait for clk_period;
x <= "000000111011011011";  
wait for clk_period;
x <= "111111011001011011";  
wait for clk_period;
x <= "000000000101011001";  
wait for clk_period;
x <= "000000111000101010";  
wait for clk_period;
x <= "111111010110011010";  
wait for clk_period;
x <= "111111011000111101";  
wait for clk_period;
x <= "111110011000000101";  
wait for clk_period;
x <= "000000001110010110";  
wait for clk_period;
x <= "111111110100001100";  
wait for clk_period;
x <= "000001110111100101";  
wait for clk_period;
x <= "111110110011010001";  
wait for clk_period;
x <= "111111010111011001";  
wait for clk_period;
x <= "111111001000100110";  
wait for clk_period;
x <= "000000001001100101";  
wait for clk_period;
x <= "111111100101100101";  
wait for clk_period;
x <= "111111011010111001";  
wait for clk_period;
x <= "000000100100101111";  
wait for clk_period;
x <= "000000110100100110";  
wait for clk_period;
x <= "000000001010101001";  
wait for clk_period;
x <= "000000100010000001";  
wait for clk_period;
x <= "000001001110100101";  
wait for clk_period;
x <= "111111110011110111";  
wait for clk_period;
x <= "000001010000111110";  
wait for clk_period;
x <= "111111010111100000";  
wait for clk_period;
x <= "000000111001101110";  
wait for clk_period;
x <= "000000111110101010";  
wait for clk_period;
x <= "000001110010001011";  
wait for clk_period;
x <= "111110011011100110";  
wait for clk_period;
x <= "111111101100110111";  
wait for clk_period;
x <= "000000100010001001";  
wait for clk_period;
x <= "111111110010011110";  
wait for clk_period;
x <= "000000001110001000";  
wait for clk_period;
x <= "111110111101011111";  
wait for clk_period;
x <= "000000011110010011";  
wait for clk_period;
x <= "000000111010001111";  
wait for clk_period;
x <= "111111001110111101";  
wait for clk_period;
x <= "111111011101011010";  
wait for clk_period;
x <= "000001000100100100";  
wait for clk_period;
x <= "000000111000101110";  
wait for clk_period;
x <= "111111011111010000";  
wait for clk_period;
x <= "000000100010001100";  
wait for clk_period;
x <= "000000101101001011";  
wait for clk_period;
x <= "111110111101011101";  
wait for clk_period;
x <= "000001100001101101";  
wait for clk_period;
x <= "111110111101011111";  
wait for clk_period;
x <= "000000000101010110";  
wait for clk_period;
x <= "111111011000111111";  
wait for clk_period;
x <= "111110011111110001";  
wait for clk_period;
x <= "111101110101100101";  
wait for clk_period;
x <= "000000000011111011";  
wait for clk_period;
x <= "000000100110000011";  
wait for clk_period;
x <= "111111000001110011";  
wait for clk_period;
x <= "111111010100100100";  
wait for clk_period;
x <= "111110010011110100";  
wait for clk_period;
x <= "000000000011000111";  
wait for clk_period;
x <= "111110110001011011";  
wait for clk_period;
x <= "000000001101000101";  
wait for clk_period;
x <= "000000000011010111";  
wait for clk_period;
x <= "000001001000100111";  
wait for clk_period;
x <= "111110110001011001";  
wait for clk_period;
x <= "000000000111011011";  
wait for clk_period;
x <= "000000010011110011";  
wait for clk_period;
x <= "111111110000011111";  
wait for clk_period;
x <= "111111110100010001";  
wait for clk_period;
x <= "111111111010001101";  
wait for clk_period;
x <= "000000110000001001";  
wait for clk_period;
x <= "000000101101011111";  
wait for clk_period;
x <= "000000011011101101";  
wait for clk_period;
x <= "111111000110100011";  
wait for clk_period;
x <= "111111111000011000";  
wait for clk_period;
x <= "111111111101000010";  
wait for clk_period;
x <= "000001000101111001";  
wait for clk_period;
x <= "111111111000110110";  
wait for clk_period;
x <= "000001000100000100";  
wait for clk_period;
x <= "000000111000101001";  
wait for clk_period;
x <= "000001110001010001";  
wait for clk_period;
x <= "111110111100011101";  
wait for clk_period;
x <= "111111011101100001";  
wait for clk_period;
x <= "000000001001111101";  
wait for clk_period;
x <= "111111111011001100";  
wait for clk_period;
x <= "000001011101111100";  
wait for clk_period;
x <= "000000010010001101";  
wait for clk_period;
x <= "000000001011100010";  
wait for clk_period;
x <= "000000000101011100";  
wait for clk_period;
x <= "000000011101000101";  
wait for clk_period;
x <= "111111110001100110";  
wait for clk_period;
x <= "111111100100100100";  
wait for clk_period;
x <= "000001000111010101";  
wait for clk_period;
x <= "000000101100100000";  
wait for clk_period;
x <= "111110111011111100";  
wait for clk_period;
x <= "000000010011001111";  
wait for clk_period;
x <= "000000011100010000";  
wait for clk_period;
x <= "000010001101001100";  
wait for clk_period;
x <= "111110011100000001";  
wait for clk_period;
x <= "111111001111110011";  
wait for clk_period;
x <= "111110110001101101";  
wait for clk_period;
x <= "000000000010011100";  
wait for clk_period;
x <= "111111011111111110";  
wait for clk_period;
x <= "111110010010110100";  
wait for clk_period;
x <= "000001001000100110";  
wait for clk_period;
x <= "000000001001100101";  
wait for clk_period;
x <= "111111110111100011";  
wait for clk_period;
x <= "111110000111101001";  
wait for clk_period;
x <= "111111011011001010";  
wait for clk_period;
x <= "111111011011101010";  
wait for clk_period;
x <= "000001101110100111";  
wait for clk_period;
x <= "000000100011010010";  
wait for clk_period;
x <= "000000101111001011";  
wait for clk_period;
x <= "000001011011101100";  
wait for clk_period;
x <= "000000101011000101";  
wait for clk_period;
x <= "111110000101010001";  
wait for clk_period;
x <= "111111110101110100";  
wait for clk_period;
x <= "000000111010111000";  
wait for clk_period;
x <= "111110111010101101";  
wait for clk_period;
x <= "000000110111010111";  
wait for clk_period;
x <= "000000011100100110";  
wait for clk_period;
x <= "111111111010111010";  
wait for clk_period;
x <= "111111100101110010";  
wait for clk_period;
x <= "111111000001011100";  
wait for clk_period;
x <= "111101111110011011";  
wait for clk_period;
x <= "111111010110000011";  
wait for clk_period;
x <= "000000010011100101";  
wait for clk_period;
x <= "000001001111110011";  
wait for clk_period;
x <= "000001000100101111";  
wait for clk_period;
x <= "000000010011100001";  
wait for clk_period;
x <= "111110100111010011";  
wait for clk_period;
x <= "000000101011100001";  
wait for clk_period;
x <= "111111111100111100";  
wait for clk_period;
x <= "111111100111101101";  
wait for clk_period;
x <= "000000100100000110";  
wait for clk_period;
x <= "111111011111111100";  
wait for clk_period;
x <= "000000100110100011";  
wait for clk_period;
x <= "000000010111110011";  
wait for clk_period;
x <= "111111100010111011";  
wait for clk_period;
x <= "111111010100110110";  
wait for clk_period;
x <= "111111101010110100";  
wait for clk_period;
x <= "111111000110111100";  
wait for clk_period;
x <= "111111000110101010";  
wait for clk_period;
x <= "111111001011000010";  
wait for clk_period;
x <= "000000110010001101";  
wait for clk_period;
x <= "000000010000111001";  
wait for clk_period;
x <= "000001101100001101";  
wait for clk_period;
x <= "111111110010000000";  
wait for clk_period;
x <= "000000110011111111";  
wait for clk_period;
x <= "111110100100101111";  
wait for clk_period;
x <= "111111001000000101";  
wait for clk_period;
x <= "000001001111010011";  
wait for clk_period;
x <= "000000000100110000";  
wait for clk_period;
x <= "000001110011001010";  
wait for clk_period;
x <= "000000101100010100";  
wait for clk_period;
x <= "000001001000011101";  
wait for clk_period;
x <= "111110100001111001";  
wait for clk_period;
x <= "000000010001000011";  
wait for clk_period;
x <= "111111101001001011";  
wait for clk_period;
x <= "000000001011100010";  
wait for clk_period;
x <= "000000101100010000";  
wait for clk_period;
x <= "000000101111011010";  
wait for clk_period;
x <= "000001110101011111";  
wait for clk_period;
x <= "000001001100000000";  
wait for clk_period;
x <= "111111110100010000";  
wait for clk_period;
x <= "111110100011111000";  
wait for clk_period;
x <= "111110111001001101";  
wait for clk_period;
x <= "111111111000010111";  
wait for clk_period;
x <= "000000111101110011";  
wait for clk_period;
x <= "000000000100010110";  
wait for clk_period;
x <= "000000000111001001";  
wait for clk_period;
x <= "111111101000010110";  
wait for clk_period;
x <= "111111101010101100";  
wait for clk_period;
x <= "111110011001011101";  
wait for clk_period;
x <= "111111000011100000";  
wait for clk_period;
x <= "000000010110000111";  
wait for clk_period;
x <= "000000010101110101";  
wait for clk_period;
x <= "111111011111001100";  
wait for clk_period;
x <= "000000111100011101";  
wait for clk_period;
x <= "111111110111110101";  
wait for clk_period;
x <= "111111011000101110";  
wait for clk_period;
x <= "111111011111110110";  
wait for clk_period;
x <= "000000100001110111";  
wait for clk_period;
x <= "111111010101101000";  
wait for clk_period;
x <= "111110111011101110";  
wait for clk_period;
x <= "000000000001010100";  
wait for clk_period;
x <= "111110110010110010";  
wait for clk_period;
x <= "111111110001000110";  
wait for clk_period;
x <= "000000010100000110";  
wait for clk_period;
x <= "111111010011001000";  
wait for clk_period;
x <= "111110110100010101";  
wait for clk_period;
x <= "111110110011100000";  
wait for clk_period;
x <= "111101110010001000";  
wait for clk_period;
x <= "000000100011010100";  
wait for clk_period;
x <= "000001000110001001";  
wait for clk_period;
x <= "000001000100001010";  
wait for clk_period;
x <= "111111111000110111";  
wait for clk_period;
x <= "000001000010110100";  
wait for clk_period;
x <= "111111111010101110";  
wait for clk_period;
x <= "000000011110111001";  
wait for clk_period;
x <= "000000001110000001";  
wait for clk_period;
x <= "111110101000000110";  
wait for clk_period;
x <= "000011010000101101";  
wait for clk_period;
x <= "000000110100110100";  
wait for clk_period;
x <= "000000111101011001";  
wait for clk_period;
x <= "111111110001011010";  
wait for clk_period;
x <= "000000011110010101";  
wait for clk_period;
x <= "111110110110001000";  
wait for clk_period;
x <= "111111000110011101";  
wait for clk_period;
x <= "000000100011110111";  
wait for clk_period;
x <= "000000011011001001";  
wait for clk_period;
x <= "000001110000111000";  
wait for clk_period;
x <= "000000011110111010";  
wait for clk_period;
x <= "111111110011011010";  
wait for clk_period;
x <= "111111110010100001";  
wait for clk_period;
x <= "111111100110101001";  
wait for clk_period;
x <= "000000001001000001";  
wait for clk_period;
x <= "000000010001010010";  
wait for clk_period;
x <= "000000101110000111";  
wait for clk_period;
x <= "000001100110101111";  
wait for clk_period;
x <= "000000010111110111";  
wait for clk_period;
x <= "111110101011011000";  
wait for clk_period;
x <= "111111001011001111";  
wait for clk_period;
x <= "000000001110101100";  
wait for clk_period;
x <= "000000000011000110";  
wait for clk_period;
x <= "000000011111100010";  
wait for clk_period;
x <= "111111000001001010";  
wait for clk_period;
x <= "111110110101000001";  
wait for clk_period;
x <= "111111101110100011";  
wait for clk_period;
x <= "000000111010001000";  
wait for clk_period;
x <= "111111010010011011";  
wait for clk_period;
x <= "111111110001001101";  
wait for clk_period;
x <= "111111110010110111";  
wait for clk_period;
x <= "111111101100100001";  
wait for clk_period;
x <= "111111111011000000";  
wait for clk_period;
x <= "111110011011010101";  
wait for clk_period;
x <= "000000010000011000";  
wait for clk_period;
x <= "000000100111111001";  
wait for clk_period;
x <= "111111011100110111";  
wait for clk_period;
x <= "111110111000100010";  
wait for clk_period;
x <= "000000010110100001";  
wait for clk_period;
x <= "111111101011000010";  
wait for clk_period;
x <= "111110110101111111";  
wait for clk_period;
x <= "111111111001111001";  
wait for clk_period;
x <= "000001000011001100";  
wait for clk_period;
x <= "000000010111011100";  
wait for clk_period;
x <= "000000101011101100";  
wait for clk_period;
x <= "111111100000111001";  
wait for clk_period;
x <= "111111101101000001";  
wait for clk_period;
x <= "000000101110000011";  
wait for clk_period;
x <= "000000000111101111";  
wait for clk_period;
x <= "000000010110110000";  
wait for clk_period;
x <= "111111101100100101";  
wait for clk_period;
x <= "000001101100010011";  
wait for clk_period;
x <= "111111011010011000";  
wait for clk_period;
x <= "111110110000011100";  
wait for clk_period;
x <= "111111100111101010";  
wait for clk_period;
x <= "111110111001000010";  
wait for clk_period;
x <= "111111110000010110";  
wait for clk_period;
x <= "111111111111101101";  
wait for clk_period;
x <= "000001100101100100";  
wait for clk_period;
x <= "000000001110000000";  
wait for clk_period;
x <= "111111011000011001";  
wait for clk_period;
x <= "111110100111101010";  
wait for clk_period;
x <= "000000000001101101";  
wait for clk_period;
x <= "000010001111110110";  
wait for clk_period;
x <= "000000000101001010";  
wait for clk_period;
x <= "000000111110101101";  
wait for clk_period;
x <= "000001000110000111";  
wait for clk_period;
x <= "111111101010101101";  
wait for clk_period;
x <= "111111011101011000";  
wait for clk_period;
x <= "111111101001011000";  
wait for clk_period;
x <= "111111011110101011";  
wait for clk_period;
x <= "000000001000101001";  
wait for clk_period;
x <= "000001000011011001";  
wait for clk_period;
x <= "111110111011011111";  
wait for clk_period;
x <= "111111001000011011";  
wait for clk_period;
x <= "000000010000111001";  
wait for clk_period;
x <= "111111101011001001";  
wait for clk_period;
x <= "111111011100110101";  
wait for clk_period;
x <= "000000101111100011";  
wait for clk_period;
x <= "000000100100000111";  
wait for clk_period;
x <= "000000101011011000";  
wait for clk_period;
x <= "000000011110001011";  
wait for clk_period;
x <= "111111101101010101";  
wait for clk_period;
x <= "000001011110100100";  
wait for clk_period;
x <= "000000111011010111";  
wait for clk_period;
x <= "000000101001011011";  
wait for clk_period;
x <= "111111101010110011";  
wait for clk_period;
x <= "111111011001001100";  
wait for clk_period;
x <= "000000111010100001";  
wait for clk_period;
x <= "000001001010101010";  
wait for clk_period;
x <= "111111011011010100";  
wait for clk_period;
x <= "111110111111000111";  
wait for clk_period;
x <= "000000111010111001";  
wait for clk_period;
x <= "000000110111110011";  
wait for clk_period;
x <= "111111000100011110";  
wait for clk_period;
x <= "111110110001000100";  
wait for clk_period;
x <= "111111001001011101";  
wait for clk_period;
x <= "000000001010011110";  
wait for clk_period;
x <= "000000101001001101";  
wait for clk_period;
x <= "111111010111111111";  
wait for clk_period;
x <= "000001001010010001";  
wait for clk_period;
x <= "000000010010011110";  
wait for clk_period;
x <= "111101110001100110";  
wait for clk_period;
x <= "111110100010000101";  
wait for clk_period;
x <= "111110101100011101";  
wait for clk_period;
x <= "000001001001111111";  
wait for clk_period;
x <= "000000101011001001";  
wait for clk_period;
x <= "000000011100010110";  
wait for clk_period;
x <= "111110010101101001";  
wait for clk_period;
x <= "000000000111010111";  
wait for clk_period;
x <= "111111101110001111";  
wait for clk_period;
x <= "111100110011110011";  
wait for clk_period;
x <= "000000110010011011";  
wait for clk_period;
x <= "000000111010111010";  
wait for clk_period;
x <= "000001011011010001";  
wait for clk_period;
x <= "000000001000010101";  
wait for clk_period;
x <= "111111100001001101";  
wait for clk_period;
x <= "111111001110110101";  
wait for clk_period;
x <= "111111010101111111";  
wait for clk_period;
x <= "000000010111111110";  
wait for clk_period;
x <= "111111010110010010";  
wait for clk_period;
x <= "000000010100110001";  
wait for clk_period;
x <= "111111111010011101";  
wait for clk_period;
x <= "111111111001110101";  
wait for clk_period;
x <= "000000011100110101";  
wait for clk_period;
x <= "000000000100110111";  
wait for clk_period;
x <= "111111101000011001";  
wait for clk_period;
x <= "111111111110000110";  
wait for clk_period;
x <= "000000011010010110";  
wait for clk_period;
x <= "000001000110010111";  
wait for clk_period;
x <= "000001001110110100";  
wait for clk_period;
x <= "000001100011110010";  
wait for clk_period;
x <= "000000110011101011";  
wait for clk_period;
x <= "000000101111001001";  
wait for clk_period;
x <= "000001010101100010";  
wait for clk_period;
x <= "000000000100110011";  
wait for clk_period;
x <= "111111111001000010";  
wait for clk_period;
x <= "000000011110101010";  
wait for clk_period;
x <= "111111001110010010";  
wait for clk_period;
x <= "111111111011101100";  
wait for clk_period;
x <= "000001011110010100";  
wait for clk_period;
x <= "000000011101100110";  
wait for clk_period;
x <= "111111001001000101";  
wait for clk_period;
x <= "111111011001000000";  
wait for clk_period;
x <= "111111000001100010";  
wait for clk_period;
x <= "111110001001100100";  
wait for clk_period;
x <= "000000010101110101";  
wait for clk_period;
x <= "000000111010010101";  
wait for clk_period;
x <= "000000111110110110";  
wait for clk_period;
x <= "000001001100001100";  
wait for clk_period;
x <= "000000100010010001";  
wait for clk_period;
x <= "111111000101111110";  
wait for clk_period;
x <= "111110110011101101";  
wait for clk_period;
x <= "111110000000010110";  
wait for clk_period;
x <= "000000110101101001";  
wait for clk_period;
x <= "000001011110010001";  
wait for clk_period;
x <= "000000110011101101";  
wait for clk_period;
x <= "111111001111100001";  
wait for clk_period;
x <= "111110101100010110";  
wait for clk_period;
x <= "111111000110111100";  
wait for clk_period;
x <= "111110001001011000";  
wait for clk_period;
x <= "111111111101011101";  
wait for clk_period;
x <= "111110100111001111";  
wait for clk_period;
x <= "000001010000100011";  
wait for clk_period;
x <= "000000000001110011";  
wait for clk_period;
x <= "111111100000010011";  
wait for clk_period;
x <= "000000010001001010";  
wait for clk_period;
x <= "111111100011100011";  
wait for clk_period;
x <= "000000011011110011";  
wait for clk_period;
x <= "111110110001101010";  
wait for clk_period;
x <= "111111111111011000";  
wait for clk_period;
x <= "000001001011001101";  
wait for clk_period;
x <= "000001011010011101";  
wait for clk_period;
x <= "111111110001010100";  
wait for clk_period;
x <= "111111110001010011";  
wait for clk_period;
x <= "000001010000011010";  
wait for clk_period;
x <= "111111011110101011";  
wait for clk_period;
x <= "111111100011010101";  
wait for clk_period;
x <= "000000101010111110";  
wait for clk_period;
x <= "111111001011111111";  
wait for clk_period;
x <= "000000101011101101";  
wait for clk_period;
x <= "000001000111000101";  
wait for clk_period;
x <= "000000010010101101";  
wait for clk_period;
x <= "000000010000011000";  
wait for clk_period;
x <= "000000110011110111";  
wait for clk_period;
x <= "111111011100000000";  
wait for clk_period;
x <= "111111101111000000";  
wait for clk_period;
x <= "111111011011100101";  
wait for clk_period;
x <= "111111001010101000";  
wait for clk_period;
x <= "000000100100100100";  
wait for clk_period;
x <= "000001101010000110";  
wait for clk_period;
x <= "000000101100101111";  
wait for clk_period;
x <= "111111010100010011";  
wait for clk_period;
x <= "111111000110110110";  
wait for clk_period;
x <= "111101111010010000";  
wait for clk_period;
x <= "000000100001101011";  
wait for clk_period;
x <= "000000011011110011";  
wait for clk_period;
x <= "000001011000010000";  
wait for clk_period;
x <= "000001110011100101";  
wait for clk_period;
x <= "000000111001101001";  
wait for clk_period;
x <= "111110101011001010";  
wait for clk_period;
x <= "111111100001011110";  
wait for clk_period;
x <= "000000110010001101";  
wait for clk_period;
x <= "000000000111000010";  
wait for clk_period;
x <= "111111100110011011";  
wait for clk_period;
x <= "000000101111001101";  
wait for clk_period;
x <= "000001001111010110";  
wait for clk_period;
x <= "111111100010101111";  
wait for clk_period;
x <= "111111110111001100";  
wait for clk_period;
x <= "111110001011110100";  
wait for clk_period;
x <= "000000000000111101";  
wait for clk_period;
x <= "111111011100001011";  
wait for clk_period;
x <= "000001010000001100";  
wait for clk_period;
x <= "111111100011110011";  
wait for clk_period;
x <= "000000010110100000";  
wait for clk_period;
x <= "000001011011101001";  
wait for clk_period;
x <= "111111111010010011";  
wait for clk_period;
x <= "000001000000011110";  
wait for clk_period;
x <= "111111010011100100";  
wait for clk_period;
x <= "000000100000100110";  
wait for clk_period;
x <= "000000100101100111";  
wait for clk_period;
x <= "000000101001010100";  
wait for clk_period;
x <= "000000001100100110";  
wait for clk_period;
x <= "111111100101010111";  
wait for clk_period;
x <= "000000001001000111";  
wait for clk_period;
x <= "111111001010001011";  
wait for clk_period;
x <= "111111011011010111";  
wait for clk_period;
x <= "111111010011100010";  
wait for clk_period;
x <= "111110001110100001";  
wait for clk_period;
x <= "111111110110110001";  
wait for clk_period;
x <= "111110001110111110";  
wait for clk_period;
x <= "111111110000010110";  
wait for clk_period;
x <= "000000101100001001";  
wait for clk_period;
x <= "000000111010111000";  
wait for clk_period;
x <= "111111000100001101";  
wait for clk_period;
x <= "111110010101011011";  
wait for clk_period;
x <= "111111011011111001";  
wait for clk_period;
x <= "000000101000111110";  
wait for clk_period;
x <= "000000010110010011";  
wait for clk_period;
x <= "111111110010101011";  
wait for clk_period;
x <= "000001000110000000";  
wait for clk_period;
x <= "111111101001100001";  
wait for clk_period;
x <= "111111011100110010";  
wait for clk_period;
x <= "111110100011111100";  
wait for clk_period;
x <= "111111101100101111";  
wait for clk_period;
x <= "111111001101101010";  
wait for clk_period;
x <= "000001111101100001";  
wait for clk_period;
x <= "111111101111000111";  
wait for clk_period;
x <= "000000001001101110";  
wait for clk_period;
x <= "000000101110101100";  
wait for clk_period;
x <= "111111001001010000";  
wait for clk_period;
x <= "111111011000000100";  
wait for clk_period;
x <= "000001001000110011";  
wait for clk_period;
x <= "000001010101110011";  
wait for clk_period;
x <= "000000000110100011";  
wait for clk_period;
x <= "000000111100110101";  
wait for clk_period;
x <= "000000000010111011";  
wait for clk_period;
x <= "000001010100100111";  
wait for clk_period;
x <= "000000000011111010";  
wait for clk_period;
x <= "111111101100001111";  
wait for clk_period;
x <= "000000000101000000";  
wait for clk_period;
x <= "000010001011001100";  
wait for clk_period;
x <= "111111100010100100";  
wait for clk_period;
x <= "000000101100101001";  
wait for clk_period;
x <= "000001011100001010";  
wait for clk_period;
x <= "111111001101110011";  
wait for clk_period;
x <= "000000010001110100";  
wait for clk_period;
x <= "000000001110110101";  
wait for clk_period;
x <= "000000101101010101";  
wait for clk_period;
x <= "000000101001000011";  
wait for clk_period;
x <= "000000001101110010";  
wait for clk_period;
x <= "111110101000111000";  
wait for clk_period;
x <= "111111000101010110";  
wait for clk_period;
x <= "000001001000111000";  
wait for clk_period;
x <= "111111101100111101";  
wait for clk_period;
x <= "111110101010001110";  
wait for clk_period;
x <= "111111100110000010";  
wait for clk_period;
x <= "111110110011101010";  
wait for clk_period;
x <= "000000000001110001";  
wait for clk_period;
x <= "111110010111111011";  
wait for clk_period;
x <= "000000010001110000";  
wait for clk_period;
x <= "111111101011111100";  
wait for clk_period;
x <= "000000100111001100";  
wait for clk_period;
x <= "111111111101110101";  
wait for clk_period;
x <= "111110100011010101";  
wait for clk_period;
x <= "111111100100101001";  
wait for clk_period;
x <= "111111110000100010";  
wait for clk_period;
x <= "000001100000111010";  
wait for clk_period;
x <= "111111110111101001";  
wait for clk_period;
x <= "000000011011101110";  
wait for clk_period;
x <= "111111001110010110";  
wait for clk_period;
x <= "111111110010100110";  
wait for clk_period;
x <= "111110001100100000";  
wait for clk_period;
x <= "111111011001111000";  
wait for clk_period;
x <= "000000001111101110";  
wait for clk_period;
x <= "000001011010110111";  
wait for clk_period;
x <= "111110100101100101";  
wait for clk_period;
x <= "111111000001011000";  
wait for clk_period;
x <= "000000010101011011";  
wait for clk_period;
x <= "000000000010010111";  
wait for clk_period;
x <= "000000000100011110";  
wait for clk_period;
x <= "111111001100101100";  
wait for clk_period;
x <= "000000111100010100";  
wait for clk_period;
x <= "000001110101110010";  
wait for clk_period;
x <= "000010010111011110";  
wait for clk_period;
x <= "111111101001000111";  
wait for clk_period;
x <= "111111101111111001";  
wait for clk_period;
x <= "000000010100110000";  
wait for clk_period;
x <= "000000111011000011";  
wait;

    end process;
    
    
    log_process : process(clk)
        file output_file : text open write_mode is "C:\Users\Francesco\Desktop\AR\_COLLABORAZIONE CON CNR\Test su Arduino\y_filtered_FPGA.txt";
        variable row  : line;
        variable y_int   : integer;
        variable counter : integer := 0;  
    begin
        if(rising_edge(clk)) then
            if rst = '0' and now >= start_time and now <= stop_time then
                y_int := to_integer(signed(y));
                write(row,  to_integer(signed(y)), left, 25);
                writeline(output_file, row);
                report "y[" & integer'image(counter) & "] = " & integer'image(y_int);            
                counter := counter + 1;
            end if;    
        end if; 
   end process;

end architecture sim;
