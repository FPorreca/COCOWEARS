library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity testbench is
--  Port ( );
end testbench;

architecture Behavioral of testbench is
    signal A1_x: std_logic_vector(7 downto 0);
    signal A1_y: std_logic_vector(7 downto 0);
    signal A2_x: std_logic_vector(7 downto 0);
    signal A2_y: std_logic_vector(7 downto 0);
    signal A3_x: std_logic_vector(7 downto 0);
    signal A3_y: std_logic_vector(7 downto 0);
    
    signal dist_1 : std_logic_vector(7 downto 0);
    signal dist_2 : std_logic_vector(7 downto 0);
    signal dist_3 : std_logic_vector(7 downto 0);
    signal clk : std_logic := '0';
    signal gen_rst : std_logic := '1';
    signal X_coord : std_logic_vector(12 downto 0);    
    signal Y_coord : std_logic_vector(12 downto 0); 
    signal writeFile_enable : std_logic := '0';
    
    constant clk_period : time := 5 ns;
    constant start_offset : Time := 347 ns;
    
    component Trilateration is
        Port ( 
            dist_1 : in STD_LOGIC_VECTOR (7 downto 0);
            dist_2 : in STD_LOGIC_VECTOR (7 downto 0);
            dist_3 : in STD_LOGIC_VECTOR (7 downto 0);
            A1_x : in STD_LOGIC_VECTOR (7 downto 0);
            A1_y : in STD_LOGIC_VECTOR (7 downto 0);
            A2_x : in STD_LOGIC_VECTOR (7 downto 0);
            A2_y : in STD_LOGIC_VECTOR (7 downto 0);
            A3_x : in STD_LOGIC_VECTOR (7 downto 0);
            A3_y : in STD_LOGIC_VECTOR (7 downto 0);
            clk : in STD_LOGIC;
            gen_rst : in STD_LOGIC;
            X_coord : out STD_LOGIC_VECTOR (12 downto 0);
            Y_coord : out STD_LOGIC_VECTOR (12 downto 0)
        );
    end component;

begin
     uut: Trilateration
        port map (
            dist_1 => dist_1,
            dist_2 => dist_2,
            dist_3 => dist_3,
            A1_x => A1_x,
            A1_y => A1_y,
            A2_x => A2_x,
            A2_y => A2_y,
            A3_x => A3_x,
            A3_y => A3_y,
            clk => clk,
            gen_rst => gen_rst,
            X_coord => X_coord, 
            Y_coord => Y_coord
        );
    
    clk_process : process
        begin
            clk <= '0';
            wait for clk_period/2;  --for 0.5 ns signal is '0'.
            clk <= '1';
            wait for clk_period/2;  --for next 0.5 ns signal is '1'.
    end process;

    stimulus: process
        begin			
		--stimulus
		wait for start_offset;		
		 A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00101011";	 -- 2.6875
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01101101";	 -- 6.8125
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01110001";	 -- 7.0625
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00110100";	 -- 3.25
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01110001";	 -- 7.0625
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01111001";	 -- 7.5625
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00110100";	 -- 3.25
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01110001";	 -- 7.0625
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01111001";	 -- 7.5625
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00101011";	 -- 2.6875
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01101101";	 -- 6.8125
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01110001";	 -- 7.0625
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00100010";	 -- 2.125
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01101010";	 -- 6.625
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01101001";	 -- 6.5625
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00011010";	 -- 1.625
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01101000";	 -- 6.5
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01100001";	 -- 6.0625
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00100010";	 -- 2.125
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01101010";	 -- 6.625
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01101001";	 -- 6.5625
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00011010";	 -- 1.625
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01101000";	 -- 6.5
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01100001";	 -- 6.0625
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00100010";	 -- 2.125
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01101010";	 -- 6.625
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01101001";	 -- 6.5625
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00100111";	 -- 2.4375
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01110011";	 -- 7.1875
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01101110";	 -- 6.875
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00101111";	 -- 2.9375
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01110110";	 -- 7.375
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01110110";	 -- 7.375
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00101011";	 -- 2.6875
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01101101";	 -- 6.8125
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01110001";	 -- 7.0625
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00101111";	 -- 2.9375
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01110110";	 -- 7.375
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01110110";	 -- 7.375
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00110101";	 -- 3.3125
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111111";	 -- 7.9375
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01111100";	 -- 7.75
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00111100";	 -- 3.75
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "10000011";	 -- 8.1875
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "10000011";	 -- 8.1875
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00111100";	 -- 3.75
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "10000011";	 -- 8.1875
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "10000011";	 -- 8.1875
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00110101";	 -- 3.3125
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111111";	 -- 7.9375
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01111100";	 -- 7.75
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00101111";	 -- 2.9375
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01110110";	 -- 7.375
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01110110";	 -- 7.375
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00110111";	 -- 3.4375
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111010";	 -- 7.625
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01111110";	 -- 7.875
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00101111";	 -- 2.9375
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01110110";	 -- 7.375
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01110110";	 -- 7.375
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00110101";	 -- 3.3125
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111111";	 -- 7.9375
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01111100";	 -- 7.75
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00101110";	 -- 2.875
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111100";	 -- 7.75
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01110100";	 -- 7.25
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00110101";	 -- 3.3125
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111111";	 -- 7.9375
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01111100";	 -- 7.75
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00110101";	 -- 3.3125
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111111";	 -- 7.9375
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01111100";	 -- 7.75
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00111100";	 -- 3.75
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "10000011";	 -- 8.1875
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "10000011";	 -- 8.1875
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00111100";	 -- 3.75
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "10000011";	 -- 8.1875
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "10000011";	 -- 8.1875
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00111100";	 -- 3.75
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "10000011";	 -- 8.1875
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "10000011";	 -- 8.1875
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00111100";	 -- 3.75
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "10000011";	 -- 8.1875
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "10000011";	 -- 8.1875
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00111100";	 -- 3.75
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "10000011";	 -- 8.1875
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "10000011";	 -- 8.1875
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00110101";	 -- 3.3125
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111111";	 -- 7.9375
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01111100";	 -- 7.75
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00110101";	 -- 3.3125
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111111";	 -- 7.9375
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01111100";	 -- 7.75
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00101111";	 -- 2.9375
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01110110";	 -- 7.375
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01110110";	 -- 7.375
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00110101";	 -- 3.3125
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111111";	 -- 7.9375
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01111100";	 -- 7.75
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00101110";	 -- 2.875
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111100";	 -- 7.75
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01110100";	 -- 7.25
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00101000";	 -- 2.5
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111011";	 -- 7.6875
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01101101";	 -- 6.8125
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00100100";	 -- 2.25
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111001";	 -- 7.5625
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01100111";	 -- 6.4375
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00100011";	 -- 2.1875
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111001";	 -- 7.5625
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01100001";	 -- 6.0625
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00011001";	 -- 1.5625
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01101111";	 -- 6.9375
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01011001";	 -- 5.5625
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00100011";	 -- 2.1875
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111001";	 -- 7.5625
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01100001";	 -- 6.0625
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00100100";	 -- 2.25
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111001";	 -- 7.5625
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01011100";	 -- 5.75
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00100111";	 -- 2.4375
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111010";	 -- 7.625
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01010111";	 -- 5.4375
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00101100";	 -- 2.75
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111100";	 -- 7.75
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01010011";	 -- 5.1875
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00110010";	 -- 3.125
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111110";	 -- 7.875
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01010000";	 -- 5.0
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00101100";	 -- 2.75
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111100";	 -- 7.75
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01010011";	 -- 5.1875
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00101100";	 -- 2.75
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111100";	 -- 7.75
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01010011";	 -- 5.1875
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00100111";	 -- 2.4375
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111010";	 -- 7.625
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01010111";	 -- 5.4375
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00100100";	 -- 2.25
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111001";	 -- 7.5625
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01011100";	 -- 5.75
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00100111";	 -- 2.4375
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111010";	 -- 7.625
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01010111";	 -- 5.4375
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00011111";	 -- 1.9375
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01110001";	 -- 7.0625
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01001110";	 -- 4.875
        wait for clk_period;
        A1_x <= "00000000";	 -- 0.0
        A1_y <= "00000000";	 -- 0.0
        dist_1 <= "00100111";	 -- 2.4375
        A2_x <= "01010110";	 -- 5.375
        A2_y <= "00000000";	 -- 0.0
        dist_2 <= "01111010";	 -- 7.625
        A3_x <= "00101011";	 -- 2.6875
        A3_y <= "00111000";	 -- 3.5
        dist_3 <= "01010111";	 -- 5.4375
		wait;
	end process stimulus;
	
	monitor : process(clk)
        use STD.TEXTIO.all;
        file F: TEXT open WRITE_MODE is "coords_by_FPGA.txt";
        variable row : LINE;
        
        begin
            if (writeFile_enable = '1') then
                if (rising_edge(clk)) then
                    WRITE (row, TO_BITVECTOR(X_coord), Right, 32);
                    WRITE (row, ';', Right, 1);
                    WRITE (row, TO_BITVECTOR(Y_coord), Right, 32);
                    WRITELINE (F, row);
                end if;
            end if;
    end process monitor;
    
    writeFile_enable_signal : process
        begin
            wait for 597ns;
            writeFile_enable <= '1';
            wait for 200ns;
            writeFile_enable <= '0';
            wait;
    end process writeFile_enable_signal;
                
end Behavioral;

